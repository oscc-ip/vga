module vga_ctrl(
    input wire clk,
    input wire resetn
);
    
endmodule
