`ifndef __VGA_TOP__
`define __VGA_TOP__
module vga_top(

);

endmodule
`endif
